library IEEE;
use     IEEE.std_logic_1164.all;

library PoC;
use     PoC.AXI4_Full.all;
use     PoC.AXI4Lite.all;


entity BlockDesign_top is
	port (
		signal Clock           : out std_logic;
		signal PL_Reset        : out std_logic;
		
		signal Config_m2s      : out T_AXI4Lite_Bus_M2S;
		signal Config_s2m      : in  T_AXI4Lite_Bus_S2M;
		
		signal Manager_m2s     : out T_AXI4_Bus_M2S_Vector;
		signal Manager_s2m     : in  T_AXI4_Bus_S2M_Vector;
		
		signal Subordinate_m2s : in  T_AXI4_Bus_M2S_Vector;
		signal Subordinate_s2m : out T_AXI4_Bus_S2M_Vector
	);
end entity;


architecture wrapper of BlockDesign_top is
	package AXI4_A40_D32 is new PoC.AXI4Full_Sized
		generic map (
			ADDRESS_BITS => 40,
			DATA_BITS    => 32,
			USER_BITS    => 16,
			ID_BITS      => 16
		);
		
	signal ConfigMM_m2s      : AXI4_A40_D32.Sized_M2S;
	signal ConfigMM_s2m      : AXI4_A40_D32.Sized_S2M;

	signal IRQs     : std_logic_vector(7 downto 0);

begin
	BD: entity work.BlochDesign_wrapper
		port map (
			Clock_0    => Clock,
			
			FPD_Clock  => Clock,
			LPD_Clock  => Clock,
			
			PL_IRQs    => IRQs,
			PL_Reset_0 => PL_Reset,
			
			Config_0_araddr  => ConfigMM_m2s.ARAddr,
			Config_0_arburst => ConfigMM_m2s.ARBurst,
			Config_0_arcache => ConfigMM_m2s.ARCache,
			Config_0_arid    => ConfigMM_m2s.ARID,
			Config_0_arlen   => ConfigMM_m2s.ARLen,
			Config_0_arlock  => ConfigMM_m2s.ARLock(0),
			Config_0_arprot  => ConfigMM_m2s.ARProt,
			Config_0_arqos   => ConfigMM_m2s.ARQoS,
			Config_0_arready => ConfigMM_s2m.ARReady,
			Config_0_arsize  => ConfigMM_m2s.ARSize,
			Config_0_aruser  => ConfigMM_m2s.ARUser,
			Config_0_arvalid => ConfigMM_m2s.ARValid,
			Config_0_awaddr  => ConfigMM_m2s.AWAddr,
			Config_0_awburst => ConfigMM_m2s.AWBurst,
			Config_0_awcache => ConfigMM_m2s.AWCache,
			Config_0_awid    => ConfigMM_m2s.AWID,
			Config_0_awlen   => ConfigMM_m2s.AWLen,
			Config_0_awlock  => ConfigMM_m2s.AWLock(0),
			Config_0_awprot  => ConfigMM_m2s.AWProt,
			Config_0_awqos   => ConfigMM_m2s.AWQoS,
			Config_0_awready => ConfigMM_s2m.AWReady,
			Config_0_awsize  => ConfigMM_m2s.AWSize,
			Config_0_awuser  => ConfigMM_m2s.AWUser,
			Config_0_awvalid => ConfigMM_m2s.AWValid,
			Config_0_bid     => ConfigMM_s2m.BID,
			Config_0_bready  => ConfigMM_m2s.BReady,
			Config_0_bresp   => ConfigMM_s2m.BResp,
			Config_0_bvalid  => ConfigMM_s2m.BValid,
			Config_0_rdata   => ConfigMM_s2m.RData,
			Config_0_rid     => ConfigMM_s2m.RID,
			Config_0_rlast   => ConfigMM_s2m.RLast,
			Config_0_rready  => ConfigMM_m2s.RReady,
			Config_0_rresp   => ConfigMM_s2m.RResp,
			Config_0_rvalid  => ConfigMM_s2m.RValid,
			Config_0_wdata   => ConfigMM_m2s.WData,
			Config_0_wlast   => ConfigMM_m2s.WLast,
			Config_0_wready  => ConfigMM_s2m.WReady,
			Config_0_wstrb   => ConfigMM_m2s.WStrb,
			Config_0_wvalid  => ConfigMM_m2s.WValid,
			
			Manager_0_araddr  => Manager_m2s(0).ARAddr,
			Manager_0_arburst => Manager_m2s(0).ARBurst,
			Manager_0_arcache => Manager_m2s(0).ARCache,
			Manager_0_arid    => Manager_m2s(0).ARID,
			Manager_0_arlen   => Manager_m2s(0).ARLen,
			Manager_0_arlock  => Manager_m2s(0).ARLock(0),
			Manager_0_arprot  => Manager_m2s(0).ARProt,
			Manager_0_arqos   => Manager_m2s(0).ARQoS,
			Manager_0_arready => Manager_s2m(0).ARReady,
			Manager_0_arsize  => Manager_m2s(0).ARSize,
			Manager_0_aruser  => Manager_m2s(0).ARUser,
			Manager_0_arvalid => Manager_m2s(0).ARValid,
			Manager_0_awaddr  => Manager_m2s(0).AWAddr,
			Manager_0_awburst => Manager_m2s(0).AWBurst,
			Manager_0_awcache => Manager_m2s(0).AWCache,
			Manager_0_awid    => Manager_m2s(0).AWID,
			Manager_0_awlen   => Manager_m2s(0).AWLen,
			Manager_0_awlock  => Manager_m2s(0).AWLock(0),
			Manager_0_awprot  => Manager_m2s(0).AWProt,
			Manager_0_awqos   => Manager_m2s(0).AWQoS,
			Manager_0_awready => Manager_s2m(0).AWReady,
			Manager_0_awsize  => Manager_m2s(0).AWSize,
			Manager_0_awuser  => Manager_m2s(0).AWUser,
			Manager_0_awvalid => Manager_m2s(0).AWValid,
			Manager_0_bid     => Manager_s2m(0).BID,
			Manager_0_bready  => Manager_m2s(0).BReady,
			Manager_0_bresp   => Manager_s2m(0).BResp,
			Manager_0_bvalid  => Manager_s2m(0).BValid,
			Manager_0_rdata   => Manager_s2m(0).RData,
			Manager_0_rid     => Manager_s2m(0).RID,
			Manager_0_rlast   => Manager_s2m(0).RLast,
			Manager_0_rready  => Manager_m2s(0).RReady,
			Manager_0_rresp   => Manager_s2m(0).RResp,
			Manager_0_rvalid  => Manager_s2m(0).RValid,
			Manager_0_wdata   => Manager_m2s(0).WData,
			Manager_0_wlast   => Manager_m2s(0).WLast,
			Manager_0_wready  => Manager_s2m(0).WReady,
			Manager_0_wstrb   => Manager_m2s(0).WStrb,
			Manager_0_wvalid  => Manager_m2s(0).WValid,
			
			Manager_1_araddr  => Manager_m2s(1).ARAddr,
			Manager_1_arburst => Manager_m2s(1).ARBurst,
			Manager_1_arcache => Manager_m2s(1).ARCache,
			Manager_1_arid    => Manager_m2s(1).ARID,
			Manager_1_arlen   => Manager_m2s(1).ARLen,
			Manager_1_arlock  => Manager_m2s(1).ARLock(0),
			Manager_1_arprot  => Manager_m2s(1).ARProt,
			Manager_1_arqos   => Manager_m2s(1).ARQoS,
			Manager_1_arready => Manager_s2m(1).ARReady,
			Manager_1_arsize  => Manager_m2s(1).ARSize,
			Manager_1_aruser  => Manager_m2s(1).ARUser,
			Manager_1_arvalid => Manager_m2s(1).ARValid,
			Manager_1_awaddr  => Manager_m2s(1).AWAddr,
			Manager_1_awburst => Manager_m2s(1).AWBurst,
			Manager_1_awcache => Manager_m2s(1).AWCache,
			Manager_1_awid    => Manager_m2s(1).AWID,
			Manager_1_awlen   => Manager_m2s(1).AWLen,
			Manager_1_awlock  => Manager_m2s(1).AWLock(0),
			Manager_1_awprot  => Manager_m2s(1).AWProt,
			Manager_1_awqos   => Manager_m2s(1).AWQoS,
			Manager_1_awready => Manager_s2m(1).AWReady,
			Manager_1_awsize  => Manager_m2s(1).AWSize,
			Manager_1_awuser  => Manager_m2s(1).AWUser,
			Manager_1_awvalid => Manager_m2s(1).AWValid,
			Manager_1_bid     => Manager_s2m(1).BID,
			Manager_1_bready  => Manager_m2s(1).BReady,
			Manager_1_bresp   => Manager_s2m(1).BResp,
			Manager_1_bvalid  => Manager_s2m(1).BValid,
			Manager_1_rdata   => Manager_s2m(1).RData,
			Manager_1_rid     => Manager_s2m(1).RID,
			Manager_1_rlast   => Manager_s2m(1).RLast,
			Manager_1_rready  => Manager_m2s(1).RReady,
			Manager_1_rresp   => Manager_s2m(1).RResp,
			Manager_1_rvalid  => Manager_s2m(1).RValid,
			Manager_1_wdata   => Manager_m2s(1).WData,
			Manager_1_wlast   => Manager_m2s(1).WLast,
			Manager_1_wready  => Manager_s2m(1).WReady,
			Manager_1_wstrb   => Manager_m2s(1).WStrb,
			Manager_1_wvalid  => Manager_m2s(1).WValid,
			
			Subordinate_0_araddr  => Subordinate_m2s(0).ARAddr,
			Subordinate_0_arburst => Subordinate_m2s(0).ARBurst,
			Subordinate_0_arcache => Subordinate_m2s(0).ARCache,
			Subordinate_0_arid    => Subordinate_m2s(0).ARID,
			Subordinate_0_arlen   => Subordinate_m2s(0).ARLen,
			Subordinate_0_arlock  => Subordinate_m2s(0).ARLock(0),
			Subordinate_0_arprot  => Subordinate_m2s(0).ARProt,
			Subordinate_0_arqos   => Subordinate_m2s(0).ARQoS,
			Subordinate_0_arready => Subordinate_s2m(0).ARReady,
			Subordinate_0_arsize  => Subordinate_m2s(0).ARSize,
			Subordinate_0_aruser  => Subordinate_m2s(0).ARUser(0),
			Subordinate_0_arvalid => Subordinate_m2s(0).ARValid,
			Subordinate_0_awaddr  => Subordinate_m2s(0).AWAddr,
			Subordinate_0_awburst => Subordinate_m2s(0).AWBurst,
			Subordinate_0_awcache => Subordinate_m2s(0).AWCache,
			Subordinate_0_awid    => Subordinate_m2s(0).AWID,
			Subordinate_0_awlen   => Subordinate_m2s(0).AWLen,
			Subordinate_0_awlock  => Subordinate_m2s(0).AWLock(0),
			Subordinate_0_awprot  => Subordinate_m2s(0).AWProt,
			Subordinate_0_awqos   => Subordinate_m2s(0).AWQoS,
			Subordinate_0_awready => Subordinate_s2m(0).AWReady,
			Subordinate_0_awsize  => Subordinate_m2s(0).AWSize,
			Subordinate_0_awuser  => Subordinate_m2s(0).AWUser(0),
			Subordinate_0_awvalid => Subordinate_m2s(0).AWValid,
			Subordinate_0_bid     => Subordinate_s2m(0).BID,
			Subordinate_0_bready  => Subordinate_m2s(0).BReady,
			Subordinate_0_bresp   => Subordinate_s2m(0).BResp,
			Subordinate_0_bvalid  => Subordinate_s2m(0).BValid,
			Subordinate_0_rdata   => Subordinate_s2m(0).RData,
			Subordinate_0_rid     => Subordinate_s2m(0).RID,
			Subordinate_0_rlast   => Subordinate_s2m(0).RLast,
			Subordinate_0_rready  => Subordinate_m2s(0).RReady,
			Subordinate_0_rresp   => Subordinate_s2m(0).RResp,
			Subordinate_0_rvalid  => Subordinate_s2m(0).RValid,
			Subordinate_0_wdata   => Subordinate_m2s(0).WData,
			Subordinate_0_wlast   => Subordinate_m2s(0).WLast,
			Subordinate_0_wready  => Subordinate_s2m(0).WReady,
			Subordinate_0_wstrb   => Subordinate_m2s(0).WStrb,
			Subordinate_0_wvalid  => Subordinate_m2s(0).WValid,

			Subordinate_1_araddr  => Subordinate_m2s(1).ARAddr,
			Subordinate_1_arburst => Subordinate_m2s(1).ARBurst,
			Subordinate_1_arcache => Subordinate_m2s(1).ARCache,
			Subordinate_1_arid    => Subordinate_m2s(1).ARID,
			Subordinate_1_arlen   => Subordinate_m2s(1).ARLen,
			Subordinate_1_arlock  => Subordinate_m2s(1).ARLock(0),
			Subordinate_1_arprot  => Subordinate_m2s(1).ARProt,
			Subordinate_1_arqos   => Subordinate_m2s(1).ARQoS,
			Subordinate_1_arready => Subordinate_s2m(1).ARReady,
			Subordinate_1_arsize  => Subordinate_m2s(1).ARSize,
			Subordinate_1_aruser  => Subordinate_m2s(1).ARUser(0),
			Subordinate_1_arvalid => Subordinate_m2s(1).ARValid,
			Subordinate_1_awaddr  => Subordinate_m2s(1).AWAddr,
			Subordinate_1_awburst => Subordinate_m2s(1).AWBurst,
			Subordinate_1_awcache => Subordinate_m2s(1).AWCache,
			Subordinate_1_awid    => Subordinate_m2s(1).AWID,
			Subordinate_1_awlen   => Subordinate_m2s(1).AWLen,
			Subordinate_1_awlock  => Subordinate_m2s(1).AWLock(0),
			Subordinate_1_awprot  => Subordinate_m2s(1).AWProt,
			Subordinate_1_awqos   => Subordinate_m2s(1).AWQoS,
			Subordinate_1_awready => Subordinate_s2m(1).AWReady,
			Subordinate_1_awsize  => Subordinate_m2s(1).AWSize,
			Subordinate_1_awuser  => Subordinate_m2s(1).AWUser(0),
			Subordinate_1_awvalid => Subordinate_m2s(1).AWValid,
			Subordinate_1_bid     => Subordinate_s2m(1).BID,
			Subordinate_1_bready  => Subordinate_m2s(1).BReady,
			Subordinate_1_bresp   => Subordinate_s2m(1).BResp,
			Subordinate_1_bvalid  => Subordinate_s2m(1).BValid,
			Subordinate_1_rdata   => Subordinate_s2m(1).RData,
			Subordinate_1_rid     => Subordinate_s2m(1).RID,
			Subordinate_1_rlast   => Subordinate_s2m(1).RLast,
			Subordinate_1_rready  => Subordinate_m2s(1).RReady,
			Subordinate_1_rresp   => Subordinate_s2m(1).RResp,
			Subordinate_1_rvalid  => Subordinate_s2m(1).RValid,
			Subordinate_1_wdata   => Subordinate_m2s(1).WData,
			Subordinate_1_wlast   => Subordinate_m2s(1).WLast,
			Subordinate_1_wready  => Subordinate_s2m(1).WReady,
			Subordinate_1_wstrb   => Subordinate_m2s(1).WStrb,
			Subordinate_1_wvalid  => Subordinate_m2s(1).WValid,

			Subordinate_2_araddr  => Subordinate_m2s(2).ARAddr,
			Subordinate_2_arburst => Subordinate_m2s(2).ARBurst,
			Subordinate_2_arcache => Subordinate_m2s(2).ARCache,
			Subordinate_2_arid    => Subordinate_m2s(2).ARID,
			Subordinate_2_arlen   => Subordinate_m2s(2).ARLen,
			Subordinate_2_arlock  => Subordinate_m2s(2).ARLock(0),
			Subordinate_2_arprot  => Subordinate_m2s(2).ARProt,
			Subordinate_2_arqos   => Subordinate_m2s(2).ARQoS,
			Subordinate_2_arready => Subordinate_s2m(2).ARReady,
			Subordinate_2_arsize  => Subordinate_m2s(2).ARSize,
			Subordinate_2_aruser  => Subordinate_m2s(2).ARUser(0),
			Subordinate_2_arvalid => Subordinate_m2s(2).ARValid,
			Subordinate_2_awaddr  => Subordinate_m2s(2).AWAddr,
			Subordinate_2_awburst => Subordinate_m2s(2).AWBurst,
			Subordinate_2_awcache => Subordinate_m2s(2).AWCache,
			Subordinate_2_awid    => Subordinate_m2s(2).AWID,
			Subordinate_2_awlen   => Subordinate_m2s(2).AWLen,
			Subordinate_2_awlock  => Subordinate_m2s(2).AWLock(0),
			Subordinate_2_awprot  => Subordinate_m2s(2).AWProt,
			Subordinate_2_awqos   => Subordinate_m2s(2).AWQoS,
			Subordinate_2_awready => Subordinate_s2m(2).AWReady,
			Subordinate_2_awsize  => Subordinate_m2s(2).AWSize,
			Subordinate_2_awuser  => Subordinate_m2s(2).AWUser(0),
			Subordinate_2_awvalid => Subordinate_m2s(2).AWValid,
			Subordinate_2_bid     => Subordinate_s2m(2).BID,
			Subordinate_2_bready  => Subordinate_m2s(2).BReady,
			Subordinate_2_bresp   => Subordinate_s2m(2).BResp,
			Subordinate_2_bvalid  => Subordinate_s2m(2).BValid,
			Subordinate_2_rdata   => Subordinate_s2m(2).RData,
			Subordinate_2_rid     => Subordinate_s2m(2).RID,
			Subordinate_2_rlast   => Subordinate_s2m(2).RLast,
			Subordinate_2_rready  => Subordinate_m2s(2).RReady,
			Subordinate_2_rresp   => Subordinate_s2m(2).RResp,
			Subordinate_2_rvalid  => Subordinate_s2m(2).RValid,
			Subordinate_2_wdata   => Subordinate_m2s(2).WData,
			Subordinate_2_wlast   => Subordinate_m2s(2).WLast,
			Subordinate_2_wready  => Subordinate_s2m(2).WReady,
			Subordinate_2_wstrb   => Subordinate_m2s(2).WStrb,
			Subordinate_2_wvalid  => Subordinate_m2s(2).WValid
		);
	
	ConvConfig : entity PoC.AXI4_to_AXI4Lite
		port map (
			Clock       => Clock,
			Reset       => PL_Reset,
			-- IN Port
			In_M2S      => ConfigMM_m2s,
			In_S2M      => ConfigMM_s2m,
			-- OUT Port
			Out_M2S     => Config_m2s,
			Out_S2M     => Config_s2m
		);
end architecture;

library IEEE;
use     IEEE.std_logic_1164.all;

entity BlockDesign_top is
	port (
		signal Clock : out std_logic
	);
end entity;

architecture wrapper of BlockDesign_top is
	signal IRQs     : std_logic_vector(7 downto 0);
	signal PL_Reset : std_logic;
begin
	BD: entity work.BlochDesign_wrapper
		port map (
			Clock_0    => Clock,
			
			FPD_Clock  => Clock,
			LPD_Clock  => Clock,
			
			PL_IRQs    => IRQs,
			PL_Reset_0 => PL_Reset
			
--			Config_0_araddr : out STD_LOGIC_VECTOR ( 39 downto 0 );
--			Config_0_arburst : out STD_LOGIC_VECTOR ( 1 downto 0 );
--			Config_0_arcache : out STD_LOGIC_VECTOR ( 3 downto 0 );
--			Config_0_arid : out STD_LOGIC_VECTOR ( 15 downto 0 );
--			Config_0_arlen : out STD_LOGIC_VECTOR ( 7 downto 0 );
--			Config_0_arlock : out STD_LOGIC;
--			Config_0_arprot : out STD_LOGIC_VECTOR ( 2 downto 0 );
--			Config_0_arqos : out STD_LOGIC_VECTOR ( 3 downto 0 );
--			Config_0_arready : in STD_LOGIC;
--			Config_0_arsize : out STD_LOGIC_VECTOR ( 2 downto 0 );
--			Config_0_aruser : out STD_LOGIC_VECTOR ( 15 downto 0 );
--			Config_0_arvalid : out STD_LOGIC;
--			Config_0_awaddr : out STD_LOGIC_VECTOR ( 39 downto 0 );
--			Config_0_awburst : out STD_LOGIC_VECTOR ( 1 downto 0 );
--			Config_0_awcache : out STD_LOGIC_VECTOR ( 3 downto 0 );
--			Config_0_awid : out STD_LOGIC_VECTOR ( 15 downto 0 );
--			Config_0_awlen : out STD_LOGIC_VECTOR ( 7 downto 0 );
--			Config_0_awlock : out STD_LOGIC;
--			Config_0_awprot : out STD_LOGIC_VECTOR ( 2 downto 0 );
--			Config_0_awqos : out STD_LOGIC_VECTOR ( 3 downto 0 );
--			Config_0_awready : in STD_LOGIC;
--			Config_0_awsize : out STD_LOGIC_VECTOR ( 2 downto 0 );
--			Config_0_awuser : out STD_LOGIC_VECTOR ( 15 downto 0 );
--			Config_0_awvalid : out STD_LOGIC;
--			Config_0_bid : in STD_LOGIC_VECTOR ( 15 downto 0 );
--			Config_0_bready : out STD_LOGIC;
--			Config_0_bresp : in STD_LOGIC_VECTOR ( 1 downto 0 );
--			Config_0_bvalid : in STD_LOGIC;
--			Config_0_rdata : in STD_LOGIC_VECTOR ( 31 downto 0 );
--			Config_0_rid : in STD_LOGIC_VECTOR ( 15 downto 0 );
--			Config_0_rlast : in STD_LOGIC;
--			Config_0_rready : out STD_LOGIC;
--			Config_0_rresp : in STD_LOGIC_VECTOR ( 1 downto 0 );
--			Config_0_rvalid : in STD_LOGIC;
--			Config_0_wdata : out STD_LOGIC_VECTOR ( 31 downto 0 );
--			Config_0_wlast : out STD_LOGIC;
--			Config_0_wready : in STD_LOGIC;
--			Config_0_wstrb : out STD_LOGIC_VECTOR ( 3 downto 0 );
--			Config_0_wvalid : out STD_LOGIC;

--			Manager_0_araddr : out STD_LOGIC_VECTOR ( 39 downto 0 );
--			Manager_0_arburst : out STD_LOGIC_VECTOR ( 1 downto 0 );
--			Manager_0_arcache : out STD_LOGIC_VECTOR ( 3 downto 0 );
--			Manager_0_arid : out STD_LOGIC_VECTOR ( 15 downto 0 );
--			Manager_0_arlen : out STD_LOGIC_VECTOR ( 7 downto 0 );
--			Manager_0_arlock : out STD_LOGIC;
--			Manager_0_arprot : out STD_LOGIC_VECTOR ( 2 downto 0 );
--			Manager_0_arqos : out STD_LOGIC_VECTOR ( 3 downto 0 );
--			Manager_0_arready : in STD_LOGIC;
--			Manager_0_arsize : out STD_LOGIC_VECTOR ( 2 downto 0 );
--			Manager_0_aruser : out STD_LOGIC_VECTOR ( 15 downto 0 );
--			Manager_0_arvalid : out STD_LOGIC;
--			Manager_0_awaddr : out STD_LOGIC_VECTOR ( 39 downto 0 );
--			Manager_0_awburst : out STD_LOGIC_VECTOR ( 1 downto 0 );
--			Manager_0_awcache : out STD_LOGIC_VECTOR ( 3 downto 0 );
--			Manager_0_awid : out STD_LOGIC_VECTOR ( 15 downto 0 );
--			Manager_0_awlen : out STD_LOGIC_VECTOR ( 7 downto 0 );
--			Manager_0_awlock : out STD_LOGIC;
--			Manager_0_awprot : out STD_LOGIC_VECTOR ( 2 downto 0 );
--			Manager_0_awqos : out STD_LOGIC_VECTOR ( 3 downto 0 );
--			Manager_0_awready : in STD_LOGIC;
--			Manager_0_awsize : out STD_LOGIC_VECTOR ( 2 downto 0 );
--			Manager_0_awuser : out STD_LOGIC_VECTOR ( 15 downto 0 );
--			Manager_0_awvalid : out STD_LOGIC;
--			Manager_0_bid : in STD_LOGIC_VECTOR ( 15 downto 0 );
--			Manager_0_bready : out STD_LOGIC;
--			Manager_0_bresp : in STD_LOGIC_VECTOR ( 1 downto 0 );
--			Manager_0_bvalid : in STD_LOGIC;
--			Manager_0_rdata : in STD_LOGIC_VECTOR ( 127 downto 0 );
--			Manager_0_rid : in STD_LOGIC_VECTOR ( 15 downto 0 );
--			Manager_0_rlast : in STD_LOGIC;
--			Manager_0_rready : out STD_LOGIC;
--			Manager_0_rresp : in STD_LOGIC_VECTOR ( 1 downto 0 );
--			Manager_0_rvalid : in STD_LOGIC;
--			Manager_0_wdata : out STD_LOGIC_VECTOR ( 127 downto 0 );
--			Manager_0_wlast : out STD_LOGIC;
--			Manager_0_wready : in STD_LOGIC;
--			Manager_0_wstrb : out STD_LOGIC_VECTOR ( 15 downto 0 );
--			Manager_0_wvalid : out STD_LOGIC;
			
--			Manager_1_araddr : out STD_LOGIC_VECTOR ( 39 downto 0 );
--			Manager_1_arburst : out STD_LOGIC_VECTOR ( 1 downto 0 );
--			Manager_1_arcache : out STD_LOGIC_VECTOR ( 3 downto 0 );
--			Manager_1_arid : out STD_LOGIC_VECTOR ( 15 downto 0 );
--			Manager_1_arlen : out STD_LOGIC_VECTOR ( 7 downto 0 );
--			Manager_1_arlock : out STD_LOGIC;
--			Manager_1_arprot : out STD_LOGIC_VECTOR ( 2 downto 0 );
--			Manager_1_arqos : out STD_LOGIC_VECTOR ( 3 downto 0 );
--			Manager_1_arready : in STD_LOGIC;
--			Manager_1_arsize : out STD_LOGIC_VECTOR ( 2 downto 0 );
--			Manager_1_aruser : out STD_LOGIC_VECTOR ( 15 downto 0 );
--			Manager_1_arvalid : out STD_LOGIC;
--			Manager_1_awaddr : out STD_LOGIC_VECTOR ( 39 downto 0 );
--			Manager_1_awburst : out STD_LOGIC_VECTOR ( 1 downto 0 );
--			Manager_1_awcache : out STD_LOGIC_VECTOR ( 3 downto 0 );
--			Manager_1_awid : out STD_LOGIC_VECTOR ( 15 downto 0 );
--			Manager_1_awlen : out STD_LOGIC_VECTOR ( 7 downto 0 );
--			Manager_1_awlock : out STD_LOGIC;
--			Manager_1_awprot : out STD_LOGIC_VECTOR ( 2 downto 0 );
--			Manager_1_awqos : out STD_LOGIC_VECTOR ( 3 downto 0 );
--			Manager_1_awready : in STD_LOGIC;
--			Manager_1_awsize : out STD_LOGIC_VECTOR ( 2 downto 0 );
--			Manager_1_awuser : out STD_LOGIC_VECTOR ( 15 downto 0 );
--			Manager_1_awvalid : out STD_LOGIC;
--			Manager_1_bid : in STD_LOGIC_VECTOR ( 15 downto 0 );
--			Manager_1_bready : out STD_LOGIC;
--			Manager_1_bresp : in STD_LOGIC_VECTOR ( 1 downto 0 );
--			Manager_1_bvalid : in STD_LOGIC;
--			Manager_1_rdata : in STD_LOGIC_VECTOR ( 127 downto 0 );
--			Manager_1_rid : in STD_LOGIC_VECTOR ( 15 downto 0 );
--			Manager_1_rlast : in STD_LOGIC;
--			Manager_1_rready : out STD_LOGIC;
--			Manager_1_rresp : in STD_LOGIC_VECTOR ( 1 downto 0 );
--			Manager_1_rvalid : in STD_LOGIC;
--			Manager_1_wdata : out STD_LOGIC_VECTOR ( 127 downto 0 );
--			Manager_1_wlast : out STD_LOGIC;
--			Manager_1_wready : in STD_LOGIC;
--			Manager_1_wstrb : out STD_LOGIC_VECTOR ( 15 downto 0 );
--			Manager_1_wvalid : out STD_LOGIC;
			
--			Subordinate_0_araddr : in STD_LOGIC_VECTOR ( 48 downto 0 );
--			Subordinate_0_arburst : in STD_LOGIC_VECTOR ( 1 downto 0 );
--			Subordinate_0_arcache : in STD_LOGIC_VECTOR ( 3 downto 0 );
--			Subordinate_0_arid : in STD_LOGIC_VECTOR ( 5 downto 0 );
--			Subordinate_0_arlen : in STD_LOGIC_VECTOR ( 7 downto 0 );
--			Subordinate_0_arlock : in STD_LOGIC;
--			Subordinate_0_arprot : in STD_LOGIC_VECTOR ( 2 downto 0 );
--			Subordinate_0_arqos : in STD_LOGIC_VECTOR ( 3 downto 0 );
--			Subordinate_0_arready : out STD_LOGIC;
--			Subordinate_0_arsize : in STD_LOGIC_VECTOR ( 2 downto 0 );
--			Subordinate_0_aruser : in STD_LOGIC;
--			Subordinate_0_arvalid : in STD_LOGIC;
--			Subordinate_0_awaddr : in STD_LOGIC_VECTOR ( 48 downto 0 );
--			Subordinate_0_awburst : in STD_LOGIC_VECTOR ( 1 downto 0 );
--			Subordinate_0_awcache : in STD_LOGIC_VECTOR ( 3 downto 0 );
--			Subordinate_0_awid : in STD_LOGIC_VECTOR ( 5 downto 0 );
--			Subordinate_0_awlen : in STD_LOGIC_VECTOR ( 7 downto 0 );
--			Subordinate_0_awlock : in STD_LOGIC;
--			Subordinate_0_awprot : in STD_LOGIC_VECTOR ( 2 downto 0 );
--			Subordinate_0_awqos : in STD_LOGIC_VECTOR ( 3 downto 0 );
--			Subordinate_0_awready : out STD_LOGIC;
--			Subordinate_0_awsize : in STD_LOGIC_VECTOR ( 2 downto 0 );
--			Subordinate_0_awuser : in STD_LOGIC;
--			Subordinate_0_awvalid : in STD_LOGIC;
--			Subordinate_0_bid : out STD_LOGIC_VECTOR ( 5 downto 0 );
--			Subordinate_0_bready : in STD_LOGIC;
--			Subordinate_0_bresp : out STD_LOGIC_VECTOR ( 1 downto 0 );
--			Subordinate_0_bvalid : out STD_LOGIC;
--			Subordinate_0_rdata : out STD_LOGIC_VECTOR ( 127 downto 0 );
--			Subordinate_0_rid : out STD_LOGIC_VECTOR ( 5 downto 0 );
--			Subordinate_0_rlast : out STD_LOGIC;
--			Subordinate_0_rready : in STD_LOGIC;
--			Subordinate_0_rresp : out STD_LOGIC_VECTOR ( 1 downto 0 );
--			Subordinate_0_rvalid : out STD_LOGIC;
--			Subordinate_0_wdata : in STD_LOGIC_VECTOR ( 127 downto 0 );
--			Subordinate_0_wlast : in STD_LOGIC;
--			Subordinate_0_wready : out STD_LOGIC;
--			Subordinate_0_wstrb : in STD_LOGIC_VECTOR ( 15 downto 0 );
--			Subordinate_0_wvalid : in STD_LOGIC;
			
--			Subordinate_1_araddr : in STD_LOGIC_VECTOR ( 48 downto 0 );
--			Subordinate_1_arburst : in STD_LOGIC_VECTOR ( 1 downto 0 );
--			Subordinate_1_arcache : in STD_LOGIC_VECTOR ( 3 downto 0 );
--			Subordinate_1_arid : in STD_LOGIC_VECTOR ( 5 downto 0 );
--			Subordinate_1_arlen : in STD_LOGIC_VECTOR ( 7 downto 0 );
--			Subordinate_1_arlock : in STD_LOGIC;
--			Subordinate_1_arprot : in STD_LOGIC_VECTOR ( 2 downto 0 );
--			Subordinate_1_arqos : in STD_LOGIC_VECTOR ( 3 downto 0 );
--			Subordinate_1_arready : out STD_LOGIC;
--			Subordinate_1_arsize : in STD_LOGIC_VECTOR ( 2 downto 0 );
--			Subordinate_1_aruser : in STD_LOGIC;
--			Subordinate_1_arvalid : in STD_LOGIC;
--			Subordinate_1_awaddr : in STD_LOGIC_VECTOR ( 48 downto 0 );
--			Subordinate_1_awburst : in STD_LOGIC_VECTOR ( 1 downto 0 );
--			Subordinate_1_awcache : in STD_LOGIC_VECTOR ( 3 downto 0 );
--			Subordinate_1_awid : in STD_LOGIC_VECTOR ( 5 downto 0 );
--			Subordinate_1_awlen : in STD_LOGIC_VECTOR ( 7 downto 0 );
--			Subordinate_1_awlock : in STD_LOGIC;
--			Subordinate_1_awprot : in STD_LOGIC_VECTOR ( 2 downto 0 );
--			Subordinate_1_awqos : in STD_LOGIC_VECTOR ( 3 downto 0 );
--			Subordinate_1_awready : out STD_LOGIC;
--			Subordinate_1_awsize : in STD_LOGIC_VECTOR ( 2 downto 0 );
--			Subordinate_1_awuser : in STD_LOGIC;
--			Subordinate_1_awvalid : in STD_LOGIC;
--			Subordinate_1_bid : out STD_LOGIC_VECTOR ( 5 downto 0 );
--			Subordinate_1_bready : in STD_LOGIC;
--			Subordinate_1_bresp : out STD_LOGIC_VECTOR ( 1 downto 0 );
--			Subordinate_1_bvalid : out STD_LOGIC;
--			Subordinate_1_rdata : out STD_LOGIC_VECTOR ( 127 downto 0 );
--			Subordinate_1_rid : out STD_LOGIC_VECTOR ( 5 downto 0 );
--			Subordinate_1_rlast : out STD_LOGIC;
--			Subordinate_1_rready : in STD_LOGIC;
--			Subordinate_1_rresp : out STD_LOGIC_VECTOR ( 1 downto 0 );
--			Subordinate_1_rvalid : out STD_LOGIC;
--			Subordinate_1_wdata : in STD_LOGIC_VECTOR ( 127 downto 0 );
--			Subordinate_1_wlast : in STD_LOGIC;
--			Subordinate_1_wready : out STD_LOGIC;
--			Subordinate_1_wstrb : in STD_LOGIC_VECTOR ( 15 downto 0 );
--			Subordinate_1_wvalid : in STD_LOGIC;
			
--			Subordinate_2_araddr : in STD_LOGIC_VECTOR ( 48 downto 0 );
--			Subordinate_2_arburst : in STD_LOGIC_VECTOR ( 1 downto 0 );
--			Subordinate_2_arcache : in STD_LOGIC_VECTOR ( 3 downto 0 );
--			Subordinate_2_arid : in STD_LOGIC_VECTOR ( 5 downto 0 );
--			Subordinate_2_arlen : in STD_LOGIC_VECTOR ( 7 downto 0 );
--			Subordinate_2_arlock : in STD_LOGIC;
--			Subordinate_2_arprot : in STD_LOGIC_VECTOR ( 2 downto 0 );
--			Subordinate_2_arqos : in STD_LOGIC_VECTOR ( 3 downto 0 );
--			Subordinate_2_arready : out STD_LOGIC;
--			Subordinate_2_arsize : in STD_LOGIC_VECTOR ( 2 downto 0 );
--			Subordinate_2_aruser : in STD_LOGIC;
--			Subordinate_2_arvalid : in STD_LOGIC;
--			Subordinate_2_awaddr : in STD_LOGIC_VECTOR ( 48 downto 0 );
--			Subordinate_2_awburst : in STD_LOGIC_VECTOR ( 1 downto 0 );
--			Subordinate_2_awcache : in STD_LOGIC_VECTOR ( 3 downto 0 );
--			Subordinate_2_awid : in STD_LOGIC_VECTOR ( 5 downto 0 );
--			Subordinate_2_awlen : in STD_LOGIC_VECTOR ( 7 downto 0 );
--			Subordinate_2_awlock : in STD_LOGIC;
--			Subordinate_2_awprot : in STD_LOGIC_VECTOR ( 2 downto 0 );
--			Subordinate_2_awqos : in STD_LOGIC_VECTOR ( 3 downto 0 );
--			Subordinate_2_awready : out STD_LOGIC;
--			Subordinate_2_awsize : in STD_LOGIC_VECTOR ( 2 downto 0 );
--			Subordinate_2_awuser : in STD_LOGIC;
--			Subordinate_2_awvalid : in STD_LOGIC;
--			Subordinate_2_bid : out STD_LOGIC_VECTOR ( 5 downto 0 );
--			Subordinate_2_bready : in STD_LOGIC;
--			Subordinate_2_bresp : out STD_LOGIC_VECTOR ( 1 downto 0 );
--			Subordinate_2_bvalid : out STD_LOGIC;
--			Subordinate_2_rdata : out STD_LOGIC_VECTOR ( 127 downto 0 );
--			Subordinate_2_rid : out STD_LOGIC_VECTOR ( 5 downto 0 );
--			Subordinate_2_rlast : out STD_LOGIC;
--			Subordinate_2_rready : in STD_LOGIC;
--			Subordinate_2_rresp : out STD_LOGIC_VECTOR ( 1 downto 0 );
--			Subordinate_2_rvalid : out STD_LOGIC;
--			Subordinate_2_wdata : in STD_LOGIC_VECTOR ( 127 downto 0 );
--			Subordinate_2_wlast : in STD_LOGIC;
--			Subordinate_2_wready : out STD_LOGIC;
--			Subordinate_2_wstrb : in STD_LOGIC_VECTOR ( 15 downto 0 );
--			Subordinate_2_wvalid : in std_logic
		);
	
end architecture;

library IEEE;
use     IEEE.std_logic_1164.all;
use     IEEE.numeric_std.all;

library Interfaces;
use     Interfaces.Axi4Common.all;
use     Interfaces.Axi4.all;
use     Interfaces.Axi4Lite.all;

library PoC;
use     PoC.AXI4_Full.all;
use     PoC.AXI4Lite.all;


entity BlockDesign_top is
	port (
		signal Clock           : out  std_logic;
		signal PL_Reset        : out  std_logic;
		
		signal Config          : view Axi4Lite_ManagerView;
		signal Managers        : view (Axi4_ManagerView)     of Axi4_Interface_Vector;
		signal Subordinates    : view (Axi4_SubordinateView) of Axi4_Interface_Vector
	);
end entity;


architecture wrapper of BlockDesign_top is
	package AXI4_A40_D32 is new Interfaces.AXI4_Generic
		generic map (
			ADDRESS_BITS => 40,
			DATA_BITS    => 32,
			USER_BITS    => 16,
			ID_BITS      => 16
		);
		
	signal ConfigMM : AXI4_A40_D32.Axi4_SizedInterface;

	signal IRQs     : std_logic_vector(7 downto 0);

begin
	BD: entity work.BlochDesign_wrapper
		port map (
			Clock_0    => Clock,
			
			FPD_Clock  => Clock,
			LPD_Clock  => Clock,
			
			PL_IRQs    => IRQs,
			PL_Reset_0 => PL_Reset,
			
			Address_Type(    Config_0_araddr)  =>                  ConfigMM.ReadAddress.Address,
			Burst_Type(      Config_0_arburst) =>                  ConfigMM.ReadAddress.Burst,
			Cache_Type(      Config_0_arcache) =>                  ConfigMM.ReadAddress.Cache,
			ID_Type(         Config_0_arid)    =>                  ConfigMM.ReadAddress.ID,
			Length_Type(     Config_0_arlen)   =>                  ConfigMM.ReadAddress.Length,
			                 Config_0_arlock   =>                  ConfigMM.ReadAddress.Lock(0),
			Protect_Type(    Config_0_arprot)  =>                  ConfigMM.ReadAddress.Protect,
			QoS_Type(        Config_0_arqos)   =>                  ConfigMM.ReadAddress.QoS,
			                 Config_0_arready  =>                  ConfigMM.ReadAddress.Ready,
			Size_Type(       Config_0_arsize)  =>                  ConfigMM.ReadAddress.Size,
			User_Type(       Config_0_aruser)  =>                  ConfigMM.ReadAddress.User,
			                 Config_0_arvalid  =>                  ConfigMM.ReadAddress.Valid,
			Address_Type(    Config_0_awaddr)  =>                  ConfigMM.WriteAddress.Address,
			Burst_Type(      Config_0_awburst) =>                  ConfigMM.WriteAddress.Burst,
			Cache_Type(      Config_0_awcache) =>                  ConfigMM.WriteAddress.Cache,
			ID_Type(         Config_0_awid)    =>                  ConfigMM.WriteAddress.ID,
			Length_Type(     Config_0_awlen)   =>                  ConfigMM.WriteAddress.Length,
			                 Config_0_awlock   =>                  ConfigMM.WriteAddress.Lock(0),
			Protect_Type(    Config_0_awprot)  =>                  ConfigMM.WriteAddress.Protect,
			QoS_Type(        Config_0_awqos)   =>                  ConfigMM.WriteAddress.QoS,
			                 Config_0_awready  =>                  ConfigMM.WriteAddress.Ready,
			Size_Type(       Config_0_awsize)  =>                  ConfigMM.WriteAddress.Size,
			User_Type(       Config_0_awuser)  =>                  ConfigMM.WriteAddress.User,
			                 Config_0_awvalid  =>                  ConfigMM.WriteAddress.Valid,
			                 Config_0_bid      => std_logic_vector(ConfigMM.WriteResponse.ID),
			                 Config_0_bready   =>                  ConfigMM.WriteResponse.Ready,
			                 Config_0_bresp    => std_logic_vector(ConfigMM.WriteResponse.Response),
			                 Config_0_bvalid   =>                  ConfigMM.WriteResponse.Valid,
			                 Config_0_rdata    => std_logic_vector(ConfigMM.ReadData.Data),
			                 Config_0_rid      => std_logic_vector(ConfigMM.ReadData.ID),
			                 Config_0_rlast    =>                  ConfigMM.ReadData.Last,
			                 Config_0_rready   =>                  ConfigMM.ReadData.Ready,
			                 Config_0_rresp    => std_logic_vector(ConfigMM.ReadData.Response),
			                 Config_0_rvalid   =>                  ConfigMM.ReadData.Valid,
			std_logic_vector(Config_0_wdata)   =>                  ConfigMM.WriteData.Data,
			                 Config_0_wlast    =>                  ConfigMM.WriteData.Last,
			                 Config_0_wready   =>                  ConfigMM.WriteData.Ready,
			Strobe_Type(     Config_0_wstrb)   =>                  ConfigMM.WriteData.Strobe,
			                 Config_0_wvalid   =>                  ConfigMM.WriteData.Valid,
			
			Address_Type(    Manager_0_araddr)  =>                  Managers(0).ReadAddress.Address,
			Burst_Type(      Manager_0_arburst) =>                  Managers(0).ReadAddress.Burst,
			Cache_Type(      Manager_0_arcache) =>                  Managers(0).ReadAddress.Cache,
			ID_Type(         Manager_0_arid)    =>                  Managers(0).ReadAddress.ID,
			Length_Type(     Manager_0_arlen)   =>                  Managers(0).ReadAddress.Length,
			                 Manager_0_arlock   =>                  Managers(0).ReadAddress.Lock(0),
			Protect_Type(    Manager_0_arprot)  =>                  Managers(0).ReadAddress.Protect,
			QoS_Type(        Manager_0_arqos)   =>                  Managers(0).ReadAddress.QoS,
			                 Manager_0_arready  =>                  Managers(0).ReadAddress.Ready,
			Size_Type(       Manager_0_arsize)  =>                  Managers(0).ReadAddress.Size,
			User_Type(       Manager_0_aruser)  =>                  Managers(0).ReadAddress.User,
			                 Manager_0_arvalid  =>                  Managers(0).ReadAddress.Valid,
			Address_Type(    Manager_0_awaddr)  =>                  Managers(0).WriteAddress.Address,
			Burst_Type(      Manager_0_awburst) =>                  Managers(0).WriteAddress.Burst,
			Cache_Type(      Manager_0_awcache) =>                  Managers(0).WriteAddress.Cache,
			ID_Type(         Manager_0_awid)    =>                  Managers(0).WriteAddress.ID,
			Length_Type(     Manager_0_awlen)   =>                  Managers(0).WriteAddress.Length,
			                 Manager_0_awlock   =>                  Managers(0).WriteAddress.Lock(0),
			Protect_Type(    Manager_0_awprot)  =>                  Managers(0).WriteAddress.Protect,
			QoS_Type(        Manager_0_awqos)   =>                  Managers(0).WriteAddress.QoS,
			                 Manager_0_awready  =>                  Managers(0).WriteAddress.Ready,
			Size_Type(       Manager_0_awsize)  =>                  Managers(0).WriteAddress.Size,
			User_Type(       Manager_0_awuser)  =>                  Managers(0).WriteAddress.User,
			                 Manager_0_awvalid  =>                  Managers(0).WriteAddress.Valid,
			                 Manager_0_bid      => std_logic_vector(Managers(0).WriteResponse.ID),
			                 Manager_0_bready   =>                  Managers(0).WriteResponse.Ready,
			                 Manager_0_bresp    => std_logic_vector(Managers(0).WriteResponse.Response),
			                 Manager_0_bvalid   =>                  Managers(0).WriteResponse.Valid,
			                 Manager_0_rdata    => std_logic_vector(Managers(0).ReadData.Data),
			                 Manager_0_rid      => std_logic_vector(Managers(0).ReadData.ID),
			                 Manager_0_rlast    =>                  Managers(0).ReadData.Last,
			                 Manager_0_rready   =>                  Managers(0).ReadData.Ready,
			                 Manager_0_rresp    => std_logic_vector(Managers(0).ReadData.Response),
			                 Manager_0_rvalid   =>                  Managers(0).ReadData.Valid,
			std_logic_vector(Manager_0_wdata)   =>                  Managers(0).WriteData.Data,
			                 Manager_0_wlast    =>                  Managers(0).WriteData.Last,
			                 Manager_0_wready   =>                  Managers(0).WriteData.Ready,
			Strobe_Type(     Manager_0_wstrb)   =>                  Managers(0).WriteData.Strobe,
			                 Manager_0_wvalid   =>                  Managers(0).WriteData.Valid,
			
			Address_Type(    Manager_1_araddr)  =>                  Managers(1).ReadAddress.Address,
			Burst_Type(      Manager_1_arburst) =>                  Managers(1).ReadAddress.Burst,
			Cache_Type(      Manager_1_arcache) =>                  Managers(1).ReadAddress.Cache,
			ID_Type(         Manager_1_arid)    =>                  Managers(1).ReadAddress.ID,
			Length_Type(     Manager_1_arlen)   =>                  Managers(1).ReadAddress.Length,
			                 Manager_1_arlock   =>                  Managers(1).ReadAddress.Lock(0),
			Protect_Type(    Manager_1_arprot)  =>                  Managers(1).ReadAddress.Protect,
			QoS_Type(        Manager_1_arqos)   =>                  Managers(1).ReadAddress.QoS,
			                 Manager_1_arready  =>                  Managers(1).ReadAddress.Ready,
			Size_Type(       Manager_1_arsize)  =>                  Managers(1).ReadAddress.Size,
			User_Type(       Manager_1_aruser)  =>                  Managers(1).ReadAddress.User,
			                 Manager_1_arvalid  =>                  Managers(1).ReadAddress.Valid,
			Address_Type(    Manager_1_awaddr)  =>                  Managers(1).WriteAddress.Address,
			Burst_Type(      Manager_1_awburst) =>                  Managers(1).WriteAddress.Burst,
			Cache_Type(      Manager_1_awcache) =>                  Managers(1).WriteAddress.Cache,
			ID_Type(         Manager_1_awid)    =>                  Managers(1).WriteAddress.ID,
			Length_Type(     Manager_1_awlen)   =>                  Managers(1).WriteAddress.Length,
			                 Manager_1_awlock   =>                  Managers(1).WriteAddress.Lock(0),
			Protect_Type(    Manager_1_awprot)  =>                  Managers(1).WriteAddress.Protect,
			QoS_Type(        Manager_1_awqos)   =>                  Managers(1).WriteAddress.QoS,
			                 Manager_1_awready  =>                  Managers(1).WriteAddress.Ready,
			Size_Type(       Manager_1_awsize)  =>                  Managers(1).WriteAddress.Size,
			User_Type(       Manager_1_awuser)  =>                  Managers(1).WriteAddress.User,
			                 Manager_1_awvalid  =>                  Managers(1).WriteAddress.Valid,
			                 Manager_1_bid      => std_logic_vector(Managers(1).WriteResponse.ID),
			                 Manager_1_bready   =>                  Managers(1).WriteResponse.Ready,
			                 Manager_1_bresp    => std_logic_vector(Managers(1).WriteResponse.Response),
			                 Manager_1_bvalid   =>                  Managers(1).WriteResponse.Valid,
			                 Manager_1_rdata    => std_logic_vector(Managers(1).ReadData.Data),
			                 Manager_1_rid      => std_logic_vector(Managers(1).ReadData.ID),
			                 Manager_1_rlast    =>                  Managers(1).ReadData.Last,
			                 Manager_1_rready   =>                  Managers(1).ReadData.Ready,
			                 Manager_1_rresp    => std_logic_vector(Managers(1).ReadData.Response),
			                 Manager_1_rvalid   =>                  Managers(1).ReadData.Valid,
			std_logic_vector(Manager_1_wdata)   =>                  Managers(1).WriteData.Data,
			                 Manager_1_wlast    =>                  Managers(1).WriteData.Last,
			                 Manager_1_wready   =>                  Managers(1).WriteData.Ready,
			Strobe_Type(     Manager_1_wstrb)   =>                  Managers(1).WriteData.Strobe,
			                 Manager_1_wvalid   =>                  Managers(1).WriteData.Valid,
			
			                 Subordinate_0_araddr   => std_logic_vector(Subordinates(0).ReadAddress.Address),
			                 Subordinate_0_arburst  => std_logic_vector(Subordinates(0).ReadAddress.Burst),
			                 Subordinate_0_arcache  => std_logic_vector(Subordinates(0).ReadAddress.Cache),
			                 Subordinate_0_arid     => std_logic_vector(Subordinates(0).ReadAddress.ID),
			                 Subordinate_0_arlen    => std_logic_vector(Subordinates(0).ReadAddress.Length),
			                 Subordinate_0_arlock   =>                  Subordinates(0).ReadAddress.Lock(0),
			                 Subordinate_0_arprot   => std_logic_vector(Subordinates(0).ReadAddress.Protect),
			                 Subordinate_0_arqos    => std_logic_vector(Subordinates(0).ReadAddress.QoS),
			                 Subordinate_0_arready  =>                  Subordinates(0).ReadAddress.Ready,
			                 Subordinate_0_arsize   => std_logic_vector(Subordinates(0).ReadAddress.Size),
			                 Subordinate_0_aruser   =>                  Subordinates(0).ReadAddress.User(0),
			                 Subordinate_0_arvalid  =>                  Subordinates(0).ReadAddress.Valid,
			                 Subordinate_0_awaddr   => std_logic_vector(Subordinates(0).WriteAddress.Address),
			                 Subordinate_0_awburst  => std_logic_vector(Subordinates(0).WriteAddress.Burst),
			                 Subordinate_0_awcache  => std_logic_vector(Subordinates(0).WriteAddress.Cache),
			                 Subordinate_0_awid     => std_logic_vector(Subordinates(0).WriteAddress.ID),
			                 Subordinate_0_awlen    => std_logic_vector(Subordinates(0).WriteAddress.Length),
			                 Subordinate_0_awlock   =>                  Subordinates(0).WriteAddress.Lock(0),
			                 Subordinate_0_awprot   => std_logic_vector(Subordinates(0).WriteAddress.Protect),
			                 Subordinate_0_awqos    => std_logic_vector(Subordinates(0).WriteAddress.QoS),
			                 Subordinate_0_awready  =>                  Subordinates(0).WriteAddress.Ready,
			                 Subordinate_0_awsize   => std_logic_vector(Subordinates(0).WriteAddress.Size),
			                 Subordinate_0_awuser   =>                  Subordinates(0).WriteAddress.User(0),
			                 Subordinate_0_awvalid  =>                  Subordinates(0).WriteAddress.Valid,
			ID_Type(         Subordinate_0_bid)     =>                  Subordinates(0).WriteResponse.ID,
			                 Subordinate_0_bready   =>                  Subordinates(0).WriteResponse.Ready,
			Response_Type(   Subordinate_0_bresp)   =>                  Subordinates(0).WriteResponse.Response,
			                 Subordinate_0_bvalid   =>                  Subordinates(0).WriteResponse.Valid,
			std_logic_vector(Subordinate_0_rdata)   =>                  Subordinates(0).ReadData.Data,
			ID_Type(         Subordinate_0_rid)     =>                  Subordinates(0).ReadData.ID,
			                 Subordinate_0_rlast    =>                  Subordinates(0).ReadData.Last,
			                 Subordinate_0_rready   =>                  Subordinates(0).ReadData.Ready,
			Response_Type(   Subordinate_0_rresp)   =>                  Subordinates(0).ReadData.Response,
			                 Subordinate_0_rvalid   =>                  Subordinates(0).ReadData.Valid,
			                 Subordinate_0_wdata    => std_logic_vector(Subordinates(0).WriteData.Data),
			                 Subordinate_0_wlast    =>                  Subordinates(0).WriteData.Last,
			                 Subordinate_0_wready   =>                  Subordinates(0).WriteData.Ready,
			                 Subordinate_0_wstrb    => std_logic_vector(Subordinates(0).WriteData.Strobe),
			                 Subordinate_0_wvalid   =>                  Subordinates(0).WriteData.Valid,
											 
			                 Subordinate_1_araddr   => std_logic_vector(Subordinates(1).ReadAddress.Address),
			                 Subordinate_1_arburst  => std_logic_vector(Subordinates(1).ReadAddress.Burst),
			                 Subordinate_1_arcache  => std_logic_vector(Subordinates(1).ReadAddress.Cache),
			                 Subordinate_1_arid     => std_logic_vector(Subordinates(1).ReadAddress.ID),
			                 Subordinate_1_arlen    => std_logic_vector(Subordinates(1).ReadAddress.Length),
			                 Subordinate_1_arlock   =>                  Subordinates(1).ReadAddress.Lock(0),
			                 Subordinate_1_arprot   => std_logic_vector(Subordinates(1).ReadAddress.Protect),
			                 Subordinate_1_arqos    => std_logic_vector(Subordinates(1).ReadAddress.QoS),
			                 Subordinate_1_arready  =>                  Subordinates(1).ReadAddress.Ready,
			                 Subordinate_1_arsize   => std_logic_vector(Subordinates(1).ReadAddress.Size),
			                 Subordinate_1_aruser   =>                  Subordinates(1).ReadAddress.User(0),
			                 Subordinate_1_arvalid  =>                  Subordinates(1).ReadAddress.Valid,
			                 Subordinate_1_awaddr   => std_logic_vector(Subordinates(1).WriteAddress.Address),
			                 Subordinate_1_awburst  => std_logic_vector(Subordinates(1).WriteAddress.Burst),
			                 Subordinate_1_awcache  => std_logic_vector(Subordinates(1).WriteAddress.Cache),
			                 Subordinate_1_awid     => std_logic_vector(Subordinates(1).WriteAddress.ID),
			                 Subordinate_1_awlen    => std_logic_vector(Subordinates(1).WriteAddress.Length),
			                 Subordinate_1_awlock   =>                  Subordinates(1).WriteAddress.Lock(0),
			                 Subordinate_1_awprot   => std_logic_vector(Subordinates(1).WriteAddress.Protect),
			                 Subordinate_1_awqos    => std_logic_vector(Subordinates(1).WriteAddress.QoS),
			                 Subordinate_1_awready  =>                  Subordinates(1).WriteAddress.Ready,
			                 Subordinate_1_awsize   => std_logic_vector(Subordinates(1).WriteAddress.Size),
			                 Subordinate_1_awuser   =>                  Subordinates(1).WriteAddress.User(0),
			                 Subordinate_1_awvalid  =>                  Subordinates(1).WriteAddress.Valid,
			ID_Type(         Subordinate_1_bid)     =>                  Subordinates(1).WriteResponse.ID,
			                 Subordinate_1_bready   =>                  Subordinates(1).WriteResponse.Ready,
			Response_Type(   Subordinate_1_bresp)   =>                  Subordinates(1).WriteResponse.Response,
			                 Subordinate_1_bvalid   =>                  Subordinates(1).WriteResponse.Valid,
			std_logic_vector(Subordinate_1_rdata)   =>                  Subordinates(1).ReadData.Data,
			ID_Type(         Subordinate_1_rid)     =>                  Subordinates(1).ReadData.ID,
			                 Subordinate_1_rlast    =>                  Subordinates(1).ReadData.Last,
			                 Subordinate_1_rready   =>                  Subordinates(1).ReadData.Ready,
			Response_Type(   Subordinate_1_rresp)   =>                  Subordinates(1).ReadData.Response,
			                 Subordinate_1_rvalid   =>                  Subordinates(1).ReadData.Valid,
			                 Subordinate_1_wdata    => std_logic_vector(Subordinates(1).WriteData.Data),
			                 Subordinate_1_wlast    =>                  Subordinates(1).WriteData.Last,
			                 Subordinate_1_wready   =>                  Subordinates(1).WriteData.Ready,
			                 Subordinate_1_wstrb    => std_logic_vector(Subordinates(1).WriteData.Strobe),
			                 Subordinate_1_wvalid   =>                  Subordinates(1).WriteData.Valid,

			                 Subordinate_2_araddr   => std_logic_vector(Subordinates(2).ReadAddress.Address),
			                 Subordinate_2_arburst  => std_logic_vector(Subordinates(2).ReadAddress.Burst),
			                 Subordinate_2_arcache  => std_logic_vector(Subordinates(2).ReadAddress.Cache),
			                 Subordinate_2_arid     => std_logic_vector(Subordinates(2).ReadAddress.ID),
			                 Subordinate_2_arlen    => std_logic_vector(Subordinates(2).ReadAddress.Length),
			                 Subordinate_2_arlock   =>                  Subordinates(2).ReadAddress.Lock(0),
			                 Subordinate_2_arprot   => std_logic_vector(Subordinates(2).ReadAddress.Protect),
			                 Subordinate_2_arqos    => std_logic_vector(Subordinates(2).ReadAddress.QoS),
			                 Subordinate_2_arready  =>                  Subordinates(2).ReadAddress.Ready,
			                 Subordinate_2_arsize   => std_logic_vector(Subordinates(2).ReadAddress.Size),
			                 Subordinate_2_aruser   =>                  Subordinates(2).ReadAddress.User(0),
			                 Subordinate_2_arvalid  =>                  Subordinates(2).ReadAddress.Valid,
			                 Subordinate_2_awaddr   => std_logic_vector(Subordinates(2).WriteAddress.Address),
			                 Subordinate_2_awburst  => std_logic_vector(Subordinates(2).WriteAddress.Burst),
			                 Subordinate_2_awcache  => std_logic_vector(Subordinates(2).WriteAddress.Cache),
			                 Subordinate_2_awid     => std_logic_vector(Subordinates(2).WriteAddress.ID),
			                 Subordinate_2_awlen    => std_logic_vector(Subordinates(2).WriteAddress.Length),
			                 Subordinate_2_awlock   =>                  Subordinates(2).WriteAddress.Lock(0),
			                 Subordinate_2_awprot   => std_logic_vector(Subordinates(2).WriteAddress.Protect),
			                 Subordinate_2_awqos    => std_logic_vector(Subordinates(2).WriteAddress.QoS),
			                 Subordinate_2_awready  =>                  Subordinates(2).WriteAddress.Ready,
			                 Subordinate_2_awsize   => std_logic_vector(Subordinates(2).WriteAddress.Size),
			                 Subordinate_2_awuser   =>                  Subordinates(2).WriteAddress.User(0),
			                 Subordinate_2_awvalid  =>                  Subordinates(2).WriteAddress.Valid,
			ID_Type(         Subordinate_2_bid)     =>                  Subordinates(2).WriteResponse.ID,
			                 Subordinate_2_bready   =>                  Subordinates(2).WriteResponse.Ready,
			Response_Type(   Subordinate_2_bresp)   =>                  Subordinates(2).WriteResponse.Response,
			                 Subordinate_2_bvalid   =>                  Subordinates(2).WriteResponse.Valid,
			std_logic_vector(Subordinate_2_rdata)   =>                  Subordinates(2).ReadData.Data,
			ID_Type(         Subordinate_2_rid)     =>                  Subordinates(2).ReadData.ID,
			                 Subordinate_2_rlast    =>                  Subordinates(2).ReadData.Last,
			                 Subordinate_2_rready   =>                  Subordinates(2).ReadData.Ready,
			Response_Type(   Subordinate_2_rresp)   =>                  Subordinates(2).ReadData.Response,
			                 Subordinate_2_rvalid   =>                  Subordinates(2).ReadData.Valid,
			                 Subordinate_2_wdata    => std_logic_vector(Subordinates(2).WriteData.Data),
			                 Subordinate_2_wlast    =>                  Subordinates(2).WriteData.Last,
			                 Subordinate_2_wready   =>                  Subordinates(2).WriteData.Ready,
			                 Subordinate_2_wstrb    => std_logic_vector(Subordinates(2).WriteData.Strobe),
			                 Subordinate_2_wvalid   =>                  Subordinates(2).WriteData.Valid
		);
	
	ConvConfig : entity PoC.AXI4_to_AXI4Lite
		port map (
			Clock       => Clock,
			Reset       => PL_Reset,
			
			Input       => ConfigMM,
			Output      => Config
		);
end architecture;
